`timescale 1ns / 1ps

module and_gate(
    input A,
    input B,
    output Y
    );
    
    assign Y = A & B;
    
endmodule